--------------------------------------------------------------------------------
-- Title : VGA Control RTL Architecture
-- Project : VGA Controller
--------------------------------------------------------------------------------
-- File : vga_ctrl_rtl.vhd
-- Author : Christoph Amon
-- Company : FH Technikum
-- Last update: 30.03.2020
-- Platform : ModelSim - Starter Edition 10.5b
--------------------------------------------------------------------------------
-- Description: VGA Control Unit
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 30.03.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

architecture rtl of vga_ctrl is

begin

end architecture rtl;
