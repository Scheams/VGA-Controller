--------------------------------------------------------------------------------
-- Title : VGA Control Entity
-- Project : VGA Controller
--------------------------------------------------------------------------------
-- File : vga_ctrl.vhd
-- Author : Christoph Amon
-- Company : FH Technikum
-- Last update: 30.03.2020
-- Platform : ModelSim - Starter Edition 10.5b
--------------------------------------------------------------------------------
-- Description: Entity for VGA Control
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 30.03.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity vga_ctrl is

  port (
    placeholder : inout std_logic
  );

end entity vga_ctrl;
