--------------------------------------------------------------------------------
-- Title : IO Control Entity
-- Project : VGA Controller
--------------------------------------------------------------------------------
-- File : io_ctrl.vhd
-- Author : Christoph Amon
-- Company : FH Technikum
-- Last update: 30.03.2020
-- Platform : ModelSim - Starter Edition 10.5b
--------------------------------------------------------------------------------
-- Description: Entity for IO Control
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 30.03.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity io_ctrl is

  port (
    placeholder : inout std_logic
  );

end entity io_ctrl;
