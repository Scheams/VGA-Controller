package pattern_gen1_pkg is



end package pattern_gen1_pkg;
