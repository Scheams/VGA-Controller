--------------------------------------------------------------------------------
-- Title : Source MUX RTL Configuration
-- Project : VGA Controller
--------------------------------------------------------------------------------
-- File : source_mux_cfg.vhd
-- Author : Christoph Amon
-- Company : FH Technikum
-- Last update: 30.03.2020
-- Platform : ModelSim - Starter Edition 10.5b
--------------------------------------------------------------------------------
-- Description: RTL configuration for Source MUX
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 30.03.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

configuration source_mux_rtl of source_mux is
  for rtl
  end for;
end configuration source_mux_rtl;
