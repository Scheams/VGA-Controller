library ieee;
use ieee.std_logic_1164.all;

entity pattern_gen1 is
  port (
    unknown : inout std_logic
  );
end entity pattern_gen1;
