architecture rtl of pattern_gen1 is

begin



end architecture rtl;
