--------------------------------------------------------------------------------
-- Title : Pattern Generator 1 RTL Configuration
-- Project : VGA Controller
--------------------------------------------------------------------------------
-- File : pattern_gen1_cfg.vhd
-- Author : Christoph Amon
-- Company : FH Technikum
-- Last update: 09.03.2020
-- Platform : ModelSim - Starter Edition 10.5b
--------------------------------------------------------------------------------
-- Description: RTL configuration for Pattern Generator 1
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 09.03.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

configuration pattern_gen1_rtl of pattern_gen1 is
  for rtl
  end for;
end configuration pattern_gen1_rtl;
