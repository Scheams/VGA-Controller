--------------------------------------------------------------------------------
-- Title :      VGA Top (Configuration)
-- Project :    VGA Controller
--------------------------------------------------------------------------------
-- File :       vga_top_cfg.vhd
-- Author :     Christoph Amon
-- Company :    FH Technikum
-- Last update: 01.04.2020
-- Platform :   ModelSim - Starter Edition 10.5b
-- Language:    VHDL 1076-2008
--------------------------------------------------------------------------------
-- Description: The "VGA Top" unit combines all elements together to one
--              VGA controller with implemented image generators.
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 01.04.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

configuration vga_top_structural of vga_top is
  for structural
  end for;
end configuration vga_top_structural;
