--------------------------------------------------------------------------------
-- Title : VGA Top Structural Architecture
-- Project : VGA Controller
--------------------------------------------------------------------------------
-- File : vga_top_structural.vhd
-- Author : Christoph Amon
-- Company : FH Technikum
-- Last update: 01.04.2020
-- Platform : ModelSim - Starter Edition 10.5b
-- Language: VHDL 1076-2008
--------------------------------------------------------------------------------
-- Description: VGA Top Unit
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 01.04.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

architecture structural of vga_top is

begin

end architecture structural;
