--------------------------------------------------------------------------------
-- Title : Pattern Generator 2 RTL Configuration
-- Project : VGA Controller
--------------------------------------------------------------------------------
-- File : pattern_gen2_cfg.vhd
-- Author : Christoph Amon
-- Company : FH Technikum
-- Last update: 29.03.2020
-- Platform : ModelSim - Starter Edition 10.5b
--------------------------------------------------------------------------------
-- Description: RTL configuration for Pattern Generator 2
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 29.03.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

configuration pattern_gen2_rtl of pattern_gen2 is
  for rtl
  end for;
end configuration pattern_gen2_rtl;
