configuration pattern_gen1_rtl of pattern_gen1 is
  for rtl
  end for;
end configuration pattern_gen1_rtl;
