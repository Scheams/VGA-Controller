--------------------------------------------------------------------------------
-- Title :      Pattern Generator 2 (Configuration)
-- Project :    VGA Controller
--------------------------------------------------------------------------------
-- File :       pattern_gen2_cfg.vhd
-- Author :     Christoph Amon
-- Company :    FH Technikum
-- Last update: 14.04.2020
-- Platform :   ModelSim - Starter Edition 10.5b, Vivado 2019.2
-- Language:    VHDL 1076-2002
--------------------------------------------------------------------------------
-- Description: The "Pattern Generator 2" unit creates a chess-like format with
--              the colours Red-Green-Blue. Over the whole frame there are
--              10 x 10 tiles.
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 29.03.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

configuration pattern_gen2_rtl of pattern_gen2 is
  for rtl
  end for;
end configuration pattern_gen2_rtl;
