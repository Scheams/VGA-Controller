--------------------------------------------------------------------------------
-- Title : IO Control RTL Configuration
-- Project : VGA Controller
--------------------------------------------------------------------------------
-- File : io_ctrl_cfg.vhd
-- Author : Christoph Amon
-- Company : FH Technikum
-- Last update: 30.03.2020
-- Platform : ModelSim - Starter Edition 10.5b
--------------------------------------------------------------------------------
-- Description: RTL configuration for IO Control
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 30.03.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

configuration io_ctrl_rtl of io_ctrl is
  for rtl
  end for;
end configuration io_ctrl_rtl;
