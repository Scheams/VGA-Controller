entity pattern_gen1_tb is
end entity pattern_gen1_tb;

architecture sim of pattern_gen1_tb is

begin



end architecture sim;
