--------------------------------------------------------------------------------
-- Title :      VGA Control (Configuration)
-- Project :    VGA Controller
--------------------------------------------------------------------------------
-- File :       vga_ctrl_cfg.vhd
-- Author :     Christoph Amon
-- Company :    FH Technikum
-- Last update: 02.04.2020
-- Platform :   ModelSim - Starter Edition 10.5b
-- Language:    VHDL 1076-2008
--------------------------------------------------------------------------------
-- Description: The "VGA Control" unit controlls the hardware operation that
--              is transfered through the VGA cable to the monitor. It takes
--              input signals like the colour information and monitor
--              specifications to perform this action.
--------------------------------------------------------------------------------
-- Revisions :
-- Date         Version  Author           Description
-- 30.03.2020   v1.0.0   Christoph Amon   Initial stage
--------------------------------------------------------------------------------

configuration vga_ctrl_rtl of vga_ctrl is
  for rtl
  end for;
end configuration vga_ctrl_rtl;
